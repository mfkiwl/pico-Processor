`timescale 1ps/1ps
module dmem(clk, reset, dmem_alu_result, dmem_in, dmem_out, dmem_write_en);

parameter d_width = 8;
parameter dmem_width = 256;

input                   clk;
input                   reset;
input                   dmem_write_en;
input  [d_width-1:0]    dmem_alu_result;
input  [d_width-1:0]    dmem_in;

output [d_width-1:0]    dmem_out;
  
wire    [d_width-1:0]    dmem_out;
reg    [d_width-1:0]    dmem_table   [dmem_width-1:0];
  

assign dmem_out = dmem_table[dmem_alu_result];

always@(posedge clk or negedge reset)
begin
	if(!reset)
	begin
	 dmem_table[0] = 0;
	 dmem_table[1] = 0;
	 dmem_table[2] = 0;
	 dmem_table[3] = 0;
	 dmem_table[4] = 0;
	 dmem_table[5] = 0;
	 dmem_table[6] = 0;
	 dmem_table[7] = 0;
	 dmem_table[8] = 0;
	 dmem_table[9] = 0;
	 dmem_table[10] = 0;
	 dmem_table[11] = 0;
	 dmem_table[12] = 0;
	 dmem_table[13] = 0;
	 dmem_table[14] = 0;
	 dmem_table[15] = 0;
	 dmem_table[16] = 0;
	 dmem_table[17] = 0;
	 dmem_table[18] = 0;
	 dmem_table[19] = 0;
	 dmem_table[20] = 0;
	 dmem_table[21] = 0;
	 dmem_table[22] = 0;
	 dmem_table[23] = 0;
	 dmem_table[24] = 0;
	 dmem_table[25] = 0;
	 dmem_table[26] = 0;
	 dmem_table[27] = 0;
	 dmem_table[28] = 0;
	 dmem_table[29] = 0;
	 dmem_table[30] = 0;
	 dmem_table[31] = 0;
	 dmem_table[32] = 0;
	 dmem_table[33] = 0;
	 dmem_table[34] = 0;
	 dmem_table[35] = 0;
	 dmem_table[36] = 0;
	 dmem_table[37] = 0;
	 dmem_table[38] = 0;
	 dmem_table[39] = 0;
	 dmem_table[40] = 0;
	 dmem_table[41] = 0;
	 dmem_table[42] = 0;
	 dmem_table[43] = 0;
	 dmem_table[44] = 0;
	 dmem_table[45] = 0;
	 dmem_table[46] = 0;
	 dmem_table[47] = 0;
	 dmem_table[48] = 0;
	 dmem_table[49] = 0;
	 dmem_table[50] = 0;
	 dmem_table[51] = 0;
	 dmem_table[52] = 0;
	 dmem_table[53] = 0;
	 dmem_table[54] = 0;
	 dmem_table[55] = 0;
	 dmem_table[56] = 0;
	 dmem_table[57] = 0;
	 dmem_table[58] = 0;
	 dmem_table[59] = 0;
	 dmem_table[60] = 0;
	 dmem_table[61] = 0;
	 dmem_table[62] = 0;
	 dmem_table[63] = 0;
	 dmem_table[64] = 0;
	 dmem_table[65] = 0;
	 dmem_table[66] = 0;
	 dmem_table[67] = 0;
	 dmem_table[68] = 0;
	 dmem_table[69] = 0;
	 dmem_table[70] = 0;
	 dmem_table[71] = 0;
	 dmem_table[72] = 0;
	 dmem_table[73] = 0;
	 dmem_table[74] = 0;
	 dmem_table[75] = 0;
	 dmem_table[76] = 0;
	 dmem_table[77] = 0;
	 dmem_table[78] = 0;
	 dmem_table[79] = 0;	
	 dmem_table[80] = 0;
	 dmem_table[81] = 0;
	 dmem_table[82] = 0;
	 dmem_table[83] = 0;
	 dmem_table[84] = 0;
	 dmem_table[85] = 0;
	 dmem_table[86] = 0;
	 dmem_table[87] = 0;
	 dmem_table[88] = 0;
	 dmem_table[89] = 0;	
	 dmem_table[90] = 0;
	 dmem_table[91] = 0;
	 dmem_table[92] = 0;
	 dmem_table[93] = 0;
	 dmem_table[94] = 0;
	 dmem_table[95] = 0;
	 dmem_table[96] = 0;
	 dmem_table[97] = 0;
	 dmem_table[98] = 0;
	 dmem_table[99] = 0;
	 dmem_table[100] = 0;
	 dmem_table[101] = 0;
	 dmem_table[102] = 0;
	 dmem_table[103] = 0;
	 dmem_table[104] = 0;
	 dmem_table[105] = 0;
	 dmem_table[106] = 0;
	 dmem_table[107] = 0;
	 dmem_table[108] = 0;
	 dmem_table[109] = 0;
	 dmem_table[110] = 0;
	 dmem_table[111] = 0;
	 dmem_table[112] = 0;
	 dmem_table[113] = 0;
	 dmem_table[114] = 0;
	 dmem_table[115] = 0;
	 dmem_table[116] = 0;
	 dmem_table[117] = 0;
	 dmem_table[118] = 0;
	 dmem_table[119] = 0;
	 dmem_table[120] = 0;
	 dmem_table[121] = 0;
	 dmem_table[122] = 0;
	 dmem_table[123] = 0;
	 dmem_table[124] = 0;
	 dmem_table[125] = 0;
	 dmem_table[126] = 0;
	 dmem_table[127] = 0;
	 dmem_table[128] = 0;
	 dmem_table[129] = 0;
	 dmem_table[130] = 0;
	 dmem_table[131] = 0;
	 dmem_table[132] = 0;
	 dmem_table[133] = 0;
	 dmem_table[134] = 0;
	 dmem_table[135] = 0;
	 dmem_table[136] = 0;
	 dmem_table[137] = 0;
	 dmem_table[138] = 0;
	 dmem_table[139] = 0;
	 dmem_table[140] = 0;
	 dmem_table[141] = 0;
	 dmem_table[142] = 0;
	 dmem_table[143] = 0;
	 dmem_table[144] = 0;
	 dmem_table[145] = 0;
	 dmem_table[146] = 0;
	 dmem_table[147] = 0;
	 dmem_table[148] = 0;
	 dmem_table[149] = 0;
	 dmem_table[150] = 0;
	 dmem_table[151] = 0;
	 dmem_table[152] = 0;
	 dmem_table[153] = 0;
	 dmem_table[154] = 0;
	 dmem_table[155] = 0;
	 dmem_table[156] = 0;
	 dmem_table[157] = 0;
	 dmem_table[158] = 0;
	 dmem_table[159] = 0;
	 dmem_table[160] = 0;
	 dmem_table[161] = 0;
	 dmem_table[162] = 0;
	 dmem_table[163] = 0;
	 dmem_table[164] = 0;
	 dmem_table[165] = 0;
	 dmem_table[166] = 0;
	 dmem_table[167] = 0;
	 dmem_table[168] = 0;
	 dmem_table[169] = 0;
	 dmem_table[170] = 0;
	 dmem_table[171] = 0;
	 dmem_table[172] = 0;
	 dmem_table[173] = 0;
	 dmem_table[174] = 0;
	 dmem_table[175] = 0;
	 dmem_table[176] = 0;
	 dmem_table[177] = 0;
	 dmem_table[178] = 0;
	 dmem_table[179] = 0;
	 dmem_table[180] = 0;
	 dmem_table[181] = 0;
	 dmem_table[182] = 0;
	 dmem_table[183] = 0;
	 dmem_table[184] = 0;
	 dmem_table[185] = 0;
	 dmem_table[186] = 0;
	 dmem_table[187] = 0;
	 dmem_table[188] = 0;
	 dmem_table[189] = 0;
	 dmem_table[190] = 0;
	 dmem_table[191] = 0;
	 dmem_table[192] = 0;
	 dmem_table[193] = 0;
	 dmem_table[194] = 0;
	 dmem_table[195] = 0;
	 dmem_table[196] = 0;
	 dmem_table[197] = 0;
	 dmem_table[198] = 0;
	 dmem_table[199] = 0;
	 dmem_table[200] = 0;
	 dmem_table[201] = 0;
	 dmem_table[202] = 0;
	 dmem_table[203] = 0;
	 dmem_table[204] = 0;
	 dmem_table[205] = 0;
	 dmem_table[206] = 0;
	 dmem_table[207] = 0;
	 dmem_table[208] = 0;
	 dmem_table[209] = 0;
	 dmem_table[210] = 0;
	 dmem_table[211] = 0;
	 dmem_table[212] = 0;
	 dmem_table[213] = 0;
	 dmem_table[214] = 0;
	 dmem_table[215] = 0;
	 dmem_table[216] = 0;
	 dmem_table[217] = 0;
	 dmem_table[218] = 0;
	 dmem_table[219] = 0;
	 dmem_table[220] = 0;
	 dmem_table[221] = 0;
	 dmem_table[222] = 0;
	 dmem_table[223] = 0;
	 dmem_table[224] = 0;
	 dmem_table[225] = 0;
	 dmem_table[226] = 0;
	 dmem_table[227] = 0;
	 dmem_table[228] = 0;
	 dmem_table[229] = 0;
	 dmem_table[230] = 0;
	 dmem_table[231] = 0;
	 dmem_table[232] = 0;
	 dmem_table[233] = 0;
	 dmem_table[234] = 0;
	 dmem_table[235] = 0;
	 dmem_table[236] = 0;
	 dmem_table[237] = 0;
	 dmem_table[238] = 0;
	 dmem_table[239] = 0;
	 dmem_table[240] = 0;
	 dmem_table[241] = 0;
	 dmem_table[242] = 0;
	 dmem_table[243] = 0;
	 dmem_table[244] = 0;
	 dmem_table[245] = 0;
	 dmem_table[246] = 0;
	 dmem_table[247] = 0;
	 dmem_table[248] = 0;
	 dmem_table[249] = 0;
	 dmem_table[250] = 0;
	 dmem_table[251] = 0;
	 dmem_table[252] = 0;
	 dmem_table[253] = 0;
	 dmem_table[254] = 0;
	 dmem_table[255] = 0;

	end
	
   else if(dmem_write_en == 1)
   begin
   dmem_table[dmem_alu_result] <= dmem_in; // STORE use alu for calculating an effective addr
   end
end
  
endmodule
